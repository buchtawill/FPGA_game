module frame10_rom(     //64 x 64 pixels
	input wire        clk,
	input wire [5:0]  col,
	input wire [5:0]  row,
	output reg [11:0] color_val
	);

	reg [5:0] colReg;
	reg [5:0] rowReg;

	always @ (posedge clk)begin
		rowReg <= row;
		colReg <= col;
	end

	always @*
	case({rowReg, colReg})
	    12'd2762: color_val = 12'd0;
	    12'd2763: color_val = 12'd0;
	    12'd2764: color_val = 12'd0;
	    12'd2765: color_val = 12'd0;
	    12'd2766: color_val = 12'd0;
	    12'd2767: color_val = 12'd0;
	    12'd2825: color_val = 12'd0;
	    12'd2826: color_val = 12'd3346;
	    12'd2827: color_val = 12'd3346;
	    12'd2828: color_val = 12'd3346;
	    12'd2829: color_val = 12'd3346;
	    12'd2830: color_val = 12'd3346;
	    12'd2831: color_val = 12'd3346;
	    12'd2832: color_val = 12'd0;
	    12'd2888: color_val = 12'd0;
	    12'd2889: color_val = 12'd3346;
	    12'd2890: color_val = 12'd3346;
	    12'd2891: color_val = 12'd3346;
	    12'd2892: color_val = 12'd3346;
	    12'd2893: color_val = 12'd3346;
	    12'd2894: color_val = 12'd3346;
	    12'd2895: color_val = 12'd3346;
	    12'd2896: color_val = 12'd3346;
	    12'd2897: color_val = 12'd0;
	    12'd2951: color_val = 12'd0;
	    12'd2952: color_val = 12'd3346;
	    12'd2953: color_val = 12'd3346;
	    12'd2954: color_val = 12'd3346;
	    12'd2955: color_val = 12'd3346;
	    12'd2956: color_val = 12'd0;
	    12'd2957: color_val = 12'd0;
	    12'd2958: color_val = 12'd0;
	    12'd2959: color_val = 12'd0;
	    12'd2960: color_val = 12'd0;
	    12'd2961: color_val = 12'd0;
	    12'd3015: color_val = 12'd0;
	    12'd3016: color_val = 12'd3346;
	    12'd3017: color_val = 12'd3346;
	    12'd3018: color_val = 12'd3346;
	    12'd3019: color_val = 12'd0;
	    12'd3020: color_val = 12'd2509;
	    12'd3021: color_val = 12'd2509;
	    12'd3026: color_val = 12'd0;
	    12'd3079: color_val = 12'd0;
	    12'd3080: color_val = 12'd3346;
	    12'd3081: color_val = 12'd3346;
	    12'd3082: color_val = 12'd0;
	    12'd3083: color_val = 12'd157;
	    12'd3084: color_val = 12'd2509;
	    12'd3085: color_val = 12'd2509;
	    12'd3086: color_val = 12'd2509;
	    12'd3090: color_val = 12'd2509;
	    12'd3091: color_val = 12'd0;
	    12'd3141: color_val = 12'd0;
	    12'd3142: color_val = 12'd0;
	    12'd3143: color_val = 12'd0;
	    12'd3144: color_val = 12'd2560;
	    12'd3145: color_val = 12'd3346;
	    12'd3146: color_val = 12'd0;
	    12'd3147: color_val = 12'd157;
	    12'd3148: color_val = 12'd2509;
	    12'd3149: color_val = 12'd2509;
	    12'd3150: color_val = 12'd2509;
	    12'd3151: color_val = 12'd2509;
	    12'd3152: color_val = 12'd2509;
	    12'd3153: color_val = 12'd2509;
	    12'd3154: color_val = 12'd2509;
	    12'd3155: color_val = 12'd0;
	    12'd3204: color_val = 12'd0;
	    12'd3205: color_val = 12'd3346;
	    12'd3206: color_val = 12'd3346;
	    12'd3207: color_val = 12'd0;
	    12'd3208: color_val = 12'd2560;
	    12'd3209: color_val = 12'd3346;
	    12'd3210: color_val = 12'd0;
	    12'd3211: color_val = 12'd157;
	    12'd3212: color_val = 12'd157;
	    12'd3213: color_val = 12'd157;
	    12'd3214: color_val = 12'd2509;
	    12'd3215: color_val = 12'd2509;
	    12'd3216: color_val = 12'd2509;
	    12'd3217: color_val = 12'd157;
	    12'd3218: color_val = 12'd157;
	    12'd3219: color_val = 12'd0;
	    12'd3268: color_val = 12'd0;
	    12'd3269: color_val = 12'd3346;
	    12'd3270: color_val = 12'd3346;
	    12'd3271: color_val = 12'd0;
	    12'd3272: color_val = 12'd2560;
	    12'd3273: color_val = 12'd3346;
	    12'd3274: color_val = 12'd3346;
	    12'd3275: color_val = 12'd0;
	    12'd3276: color_val = 12'd157;
	    12'd3277: color_val = 12'd157;
	    12'd3278: color_val = 12'd157;
	    12'd3279: color_val = 12'd157;
	    12'd3280: color_val = 12'd157;
	    12'd3281: color_val = 12'd157;
	    12'd3282: color_val = 12'd0;
	    12'd3332: color_val = 12'd0;
	    12'd3333: color_val = 12'd3346;
	    12'd3334: color_val = 12'd2560;
	    12'd3335: color_val = 12'd0;
	    12'd3336: color_val = 12'd2560;
	    12'd3337: color_val = 12'd3346;
	    12'd3338: color_val = 12'd3346;
	    12'd3339: color_val = 12'd3346;
	    12'd3340: color_val = 12'd0;
	    12'd3341: color_val = 12'd0;
	    12'd3342: color_val = 12'd0;
	    12'd3343: color_val = 12'd0;
	    12'd3344: color_val = 12'd0;
	    12'd3345: color_val = 12'd0;
	    12'd3346: color_val = 12'd0;
	    12'd3396: color_val = 12'd0;
	    12'd3397: color_val = 12'd2560;
	    12'd3398: color_val = 12'd2560;
	    12'd3399: color_val = 12'd0;
	    12'd3400: color_val = 12'd2560;
	    12'd3401: color_val = 12'd3346;
	    12'd3402: color_val = 12'd3346;
	    12'd3403: color_val = 12'd3346;
	    12'd3404: color_val = 12'd3346;
	    12'd3405: color_val = 12'd3346;
	    12'd3406: color_val = 12'd3346;
	    12'd3407: color_val = 12'd3346;
	    12'd3408: color_val = 12'd3346;
	    12'd3409: color_val = 12'd3346;
	    12'd3410: color_val = 12'd0;
	    12'd3460: color_val = 12'd0;
	    12'd3461: color_val = 12'd2560;
	    12'd3462: color_val = 12'd2560;
	    12'd3463: color_val = 12'd0;
	    12'd3464: color_val = 12'd2560;
	    12'd3465: color_val = 12'd2560;
	    12'd3466: color_val = 12'd3346;
	    12'd3467: color_val = 12'd3346;
	    12'd3468: color_val = 12'd3346;
	    12'd3469: color_val = 12'd3346;
	    12'd3470: color_val = 12'd3346;
	    12'd3471: color_val = 12'd3346;
	    12'd3472: color_val = 12'd3346;
	    12'd3473: color_val = 12'd3346;
	    12'd3474: color_val = 12'd0;
	    12'd3524: color_val = 12'd0;
	    12'd3525: color_val = 12'd2560;
	    12'd3526: color_val = 12'd2560;
	    12'd3527: color_val = 12'd0;
	    12'd3528: color_val = 12'd2560;
	    12'd3529: color_val = 12'd2560;
	    12'd3530: color_val = 12'd2560;
	    12'd3531: color_val = 12'd3346;
	    12'd3532: color_val = 12'd3346;
	    12'd3533: color_val = 12'd3346;
	    12'd3534: color_val = 12'd3346;
	    12'd3535: color_val = 12'd3346;
	    12'd3536: color_val = 12'd3346;
	    12'd3537: color_val = 12'd2560;
	    12'd3538: color_val = 12'd0;
	    12'd3588: color_val = 12'd0;
	    12'd3589: color_val = 12'd2560;
	    12'd3590: color_val = 12'd2560;
	    12'd3591: color_val = 12'd0;
	    12'd3592: color_val = 12'd2560;
	    12'd3593: color_val = 12'd2560;
	    12'd3594: color_val = 12'd2560;
	    12'd3595: color_val = 12'd3346;
	    12'd3596: color_val = 12'd3346;
	    12'd3597: color_val = 12'd3346;
	    12'd3598: color_val = 12'd3346;
	    12'd3599: color_val = 12'd3346;
	    12'd3600: color_val = 12'd2560;
	    12'd3601: color_val = 12'd2560;
	    12'd3602: color_val = 12'd0;
	    12'd3652: color_val = 12'd0;
	    12'd3653: color_val = 12'd2560;
	    12'd3654: color_val = 12'd2560;
	    12'd3655: color_val = 12'd0;
	    12'd3656: color_val = 12'd2560;
	    12'd3657: color_val = 12'd2560;
	    12'd3658: color_val = 12'd2560;
	    12'd3659: color_val = 12'd2560;
	    12'd3660: color_val = 12'd2560;
	    12'd3661: color_val = 12'd2560;
	    12'd3662: color_val = 12'd2560;
	    12'd3663: color_val = 12'd2560;
	    12'd3664: color_val = 12'd2560;
	    12'd3665: color_val = 12'd2560;
	    12'd3666: color_val = 12'd0;
	    12'd3716: color_val = 12'd0;
	    12'd3717: color_val = 12'd2560;
	    12'd3718: color_val = 12'd2560;
	    12'd3719: color_val = 12'd0;
	    12'd3720: color_val = 12'd2560;
	    12'd3721: color_val = 12'd2560;
	    12'd3722: color_val = 12'd2560;
	    12'd3723: color_val = 12'd2560;
	    12'd3724: color_val = 12'd2560;
	    12'd3725: color_val = 12'd2560;
	    12'd3726: color_val = 12'd2560;
	    12'd3727: color_val = 12'd2560;
	    12'd3728: color_val = 12'd2560;
	    12'd3729: color_val = 12'd2560;
	    12'd3730: color_val = 12'd0;
	    12'd3781: color_val = 12'd0;
	    12'd3782: color_val = 12'd0;
	    12'd3783: color_val = 12'd0;
	    12'd3784: color_val = 12'd2560;
	    12'd3785: color_val = 12'd2560;
	    12'd3786: color_val = 12'd2560;
	    12'd3787: color_val = 12'd2560;
	    12'd3788: color_val = 12'd2560;
	    12'd3789: color_val = 12'd2560;
	    12'd3790: color_val = 12'd2560;
	    12'd3791: color_val = 12'd2560;
	    12'd3792: color_val = 12'd2560;
	    12'd3793: color_val = 12'd2560;
	    12'd3794: color_val = 12'd0;
	    12'd3847: color_val = 12'd0;
	    12'd3848: color_val = 12'd2560;
	    12'd3849: color_val = 12'd2560;
	    12'd3850: color_val = 12'd2560;
	    12'd3851: color_val = 12'd0;
	    12'd3852: color_val = 12'd0;
	    12'd3853: color_val = 12'd0;
	    12'd3854: color_val = 12'd0;
	    12'd3855: color_val = 12'd2560;
	    12'd3856: color_val = 12'd2560;
	    12'd3857: color_val = 12'd2560;
	    12'd3858: color_val = 12'd0;
	    12'd3911: color_val = 12'd0;
	    12'd3912: color_val = 12'd2560;
	    12'd3913: color_val = 12'd2560;
	    12'd3914: color_val = 12'd2560;
	    12'd3915: color_val = 12'd0;
	    12'd3918: color_val = 12'd0;
	    12'd3919: color_val = 12'd2560;
	    12'd3920: color_val = 12'd2560;
	    12'd3921: color_val = 12'd2560;
	    12'd3922: color_val = 12'd0;
	    12'd3975: color_val = 12'd0;
	    12'd3976: color_val = 12'd2560;
	    12'd3977: color_val = 12'd2560;
	    12'd3978: color_val = 12'd2560;
	    12'd3979: color_val = 12'd0;
	    12'd3982: color_val = 12'd0;
	    12'd3983: color_val = 12'd2560;
	    12'd3984: color_val = 12'd2560;
	    12'd3985: color_val = 12'd2560;
	    12'd3986: color_val = 12'd0;
	    12'd4040: color_val = 12'd0;
	    12'd4041: color_val = 12'd0;
	    12'd4042: color_val = 12'd0;
	    12'd4047: color_val = 12'd0;
	    12'd4048: color_val = 12'd0;
	    12'd4049: color_val = 12'd0;

		default:  color_val = 12'b111111111111;
		endcase

endmodule //frame10_rom